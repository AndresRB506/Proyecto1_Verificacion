// tb_params.vh - (reservado para defines globales)

// tb_params.vh - Incluye de utilería (reservado para defines globales, actualmente vacío)
